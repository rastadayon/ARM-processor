`include "Constants"

module ConditionCheck (
    ports
);
    
endmodule